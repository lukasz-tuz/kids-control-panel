.title KiCad schematic
SW1 GND Net-_A1-Pad17_ TACT-SWITCH
SW2 GND Net-_A1-Pad18_ TACT-SWITCH
SW3 GND Net-_A1-Pad19_ TACT-SWITCH
SW4 GND Net-_A1-Pad20_ TACT-SWITCH
SW5 Net-_A1-Pad12_ KY-040
U1 NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 CA56-12SURKWA
U3 GND +3V3 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 NC_21 NC_22 NC_23 /I2C_SDA /I2C_SCL NC_24 NC_25 NC_26 NC_27 NC_28 GND +3V3 NC_29 NC_30 NC_31 NC_32 NC_33 NC_34 NC_35 NC_36 NC_37 NC_38 NC_39 NC_40 NC_41 NC_42 NC_43 NC_44 NC_45 NC_46 TFT LCD
96BB2-006-F1 /KPD0_OUT7 4x4_Keypad
U2 /KPD0_OUT0 /KPD0_OUT1 /KPD0_OUT2 /KPD0_OUT3 /KPD0_OUT4 /KPD0_OUT5 /KPD0_OUT6 /KPD0_OUT7 NC_47 GND NC_48 /I2C_SCL /I2C_SDA NC_49 GND GND GND Net-_A1-Pad26_ Net-_A1-Pad28_ Net-_A1-Pad27_ /KPD1_OUT0 /KPD1_OUT1 /KPD1_OUT2 /KPD1_OUT3 /KPD1_OUT4 /KPD1_OUT5 /KPD1_OUT6 /KPD1_OUT7 MCP23017_SP Expander Module
96BB2-006-F2 /KPD1_OUT7 4x4_Keypad
A1 NC_50 NC_51 NC_52 +3V3 +5V GND GND NC_53 NC_54 Net-_A1-Pad10_ Net-_A1-Pad11_ Net-_A1-Pad12_ /I2C_SDA /I2C_SCL NC_55 NC_56 Net-_A1-Pad17_ Net-_A1-Pad18_ Net-_A1-Pad19_ Net-_A1-Pad20_ NC_57 NC_58 NC_59 NC_60 NC_61 Net-_A1-Pad26_ Net-_A1-Pad27_ Net-_A1-Pad28_ GND NC_62 NC_63 NC_64 Arduino_UNO_R3
D1 GND /LED Matrix/LED_PWM LED
D2 GND /LED Matrix/LED_PWM LED
D3 GND /LED Matrix/LED_PWM LED
D4 GND /LED Matrix/LED_PWM LED
D5 GND /LED Matrix/LED_PWM LED
V1 /LED Matrix/LED_PWM GND VSOURCE
.end
